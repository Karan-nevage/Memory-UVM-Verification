// File: mem_sqr.sv
// Description: Defines the sequencer typedef for memory transactions.
// Sequencer typedef for memory transactions
//=======================================================================
typedef uvm_sequencer#(mem_tx) mem_sqr;
//=======================================================================